`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/09/2022 03:58:21 PM
// Design Name: 
// Module Name: full_1bit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: This module includes 1 bit full adder 
//              There are two half adders to add input bits and carry in bit
//              The carry out bit is generated by performing OR operation on carry out bits of both half adders        
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module full_1bit(
    input a,            //input bit a
    input b,            //input bit b
    input c_i,          //input carry in 
    output sum,         //output sum bit
    output c_o          //output carry bit
    );
    
    wire s_h, c_h,c_hi;
    
  half_add HA1(a, b, s_h, c_h);         //half adder to add input bits
  half_add HA2(s_h, c_i, sum, c_hi);    //half adder to add result of input bit addition and carry in bit
  or o1(c_o, c_h, c_hi);                // or gate to generate final carry out bit
endmodule
